// config_pkg.sv
package config_pkg;

  // 🌟 Set your alias here (max 20 characters)
  parameter string VALET_ALIAS = "InsertYourAliasHere";

  // 🔧 Optional: Set your logging style (Basic, Verbose, Theatrical)
  parameter string LOG_STYLE = "Theatrical";

  // 🎨 Optional: Choose your valet persona
  parameter string VALET_PERSONA = "Strategist";  // Options: "Strategist", "Gambler", "Minimalist", "Reckless"

endpackage
