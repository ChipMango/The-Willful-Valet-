if (match_vector.countones() > 1)
  $display("⚠️ CAM MULTI-MATCH WARNING: tag = %h", match_tag);